`include "pixel_interface.sv"
`include "ppi_interface.sv"
`include "svt_ahb_if.svi"



`include "svt_ahb.uvm.pkg"

`include "uvm_pkg.sv"

package cs_mipi_dsi_test_pkg;

import uvm_pkg::*;
import svt_uvm_pkg::*;
import svt_amba_common_uvm_pkg::*;
import svt_ahb_uvm_pkg::*;

`include "pixel_config.sv"
`include "ppi_config.sv"
`include "cust_svt_ahb_system_configuration.sv"
//`include "cs_mipi_config.sv"

`include "pixel_xtn.sv"
`include "ppi_transanction.sv"
`include "pixel_driver.sv"
`include "pixel_monitor.sv"
`include "pixel_sequencer.sv"
`include "pixel_sequence.sv"
//`include "amba_pv_master.sv"
//`include "ahb_virtual_sequencer.sv"
`include "ahb_master_random_discrete_virtual_sequence.sv"
`include "ahb_null_virtual_sequence.sv"
`include "ahb_master_directed_sequence.sv"

`include "ahb_master_random_discrete_virtual_sequence.sv"


`include "ppi_monitor.sv"

`include "ppi_agent.sv"
`include "pixel_agent.sv"
`include "ppi_env.sv"
`include "pixel_env.sv"
`include "ahb_uvc_env.sv"

`include "scoreboard.sv"

`include "cs_mipi_dsi_env.sv"
`include "cs_mipi_dsi_base_test.sv"


endpackage