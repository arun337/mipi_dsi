class dsi_reg_block;
  
  logic [31:0] payload;
  logic [31:0] dsi_cmd;
  logic [31:0] dsi_lng;
  logic [31:0] dsi_ctrl0;
  logic [31:0] dsi_ctrl1;
  logic [31:0] dsi_ctrl2;
  logic [31:0] dsi_ctrl3;
  logic [31:0] dsi_ctrl4;
  logic [31:0] dsi_ctrl5;
  logic [31:0] rx_cmd_data;
  logic [31:0] rx_cmd;
  logic [31:0] rd_cmd_wc;
  logic [31:0] rd_cmd_err;
  
endclass
