package ahb_uvc_pkg;
  import uvm_pkg::*;
  `include "uvm_macros.svh"
  import svt_ahb_uvm_pkg::*;
`include "cust_svt_ahb_system_configuration.sv"


`include "ahb_basic_wr_rd_seq.sv"

  `include "ahb_uvc_env.sv"
endpackage